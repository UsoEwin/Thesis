
// full datapath, includes: 
//	ll/ps/ne comp modules, controllers, and filters(in future)


// under testing

module datapath #(
	parameter input_width = 16, //overall 
	//for ne and sp
	parameter unit_width = 32,
	parameter mid_width = 37,
	parameter output_width = 40,
	//for ll
	parameter ll_mid_width = 22,
	parameter ll_output_width = 25
)(
	input
	
)	
	
	//filters

	//computing module

endmodule

